// -------------------------------------------------------------
//    Copyright 2025 Chad Quickstad
//    All Rights Reserved Worldwide
//
//    Licensed under the Apache License, Version 2.0 (the
//    "License"); you may not use this file except in
//    compliance with the License.  You may obtain a copy of
//    the License at
//
//        http://www.apache.org/licenses/LICENSE-2.0
//
//    Unless required by applicable law or agreed to in
//    writing, software distributed under the License is
//    distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//    CONDITIONS OF ANY KIND, either express or implied.  See
//    the License for the specific language governing
//    permissions and limitations under the License.
// -------------------------------------------------------------

`ifndef __UVM_ENUM_PKG_SV__
`define __UVM_ENUM_PKG_SV__

`include "uvm_macros.svh"

package uvm_enum_pkg;
    import uvm_pkg::*;
    `include "uvm_enum_macros.sv"
    `include "uvm_enum.sv"
    `include "uvm_rand_enum.sv"
endpackage

`endif
